interface DUT_IF(input bit Clock);
  logic ChipSelect;
  logic WriteEnable;
endinterface : DUT_IF
