// Package of parameters to be shared by DUT and Testbench
package common_pkg;
  parameter WordSize1 = 32;
  parameter WordSize2 = 16;
endpackage
