// abstract class interface
package probe_pkg;
  import uvm_pkg::*;

  `include "probe_abstract.sv"
endpackage : probe_pkg
